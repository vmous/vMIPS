----------------------------------------------------------------------------------
-- Company:        National and Kapodistrian University of Athens
-- Engineer:       Vassilis S. Moustakas
-- 
-- Create Date:    13:23:27 08/13/2009 
-- Design Name: 
-- Module Name:    IMEM_BR512X32 - IMEM_BR512X32_BEH 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description:    Instruction Memory Block RAM
--                 with "False" Synchronous Read
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity IMEM_BR512X32 is
    port(
        CLK : in STD_LOGIC;
        ADDR : in STD_LOGIC_VECTOR(8 downto 0);
        WE : in STD_LOGIC;
        DI : in STD_LOGIC_VECTOR(31 downto 0);
        DO : out STD_LOGIC_VECTOR(31 downto 0)
    );
end IMEM_BR512X32;

architecture IMEM_BR512X32_BEH of IMEM_BR512X32 is

    type br512x32_t is array(511 downto 0) of STD_LOGIC_VECTOR(31 downto 0);
    signal imem : br512x32_t := (

        ---------------------
        ----- Fibonacci -----
        ---------------------
        --0 => X"34040000",
        --1 => X"34010001",
        --2 => X"34020002", 
        --3 => X"34030005",
        --4 => X"A0840000",
        --5 => X"20840001",
        --6 => X"A0840000",
        --7 => X"20840001",
        --8 => X"808AFFFE",
        --9 => X"808BFFFF",
        --10 => X"014B6020",
        --11 => X"A08C0000",
        --12 => X"20840001",
        --13 => X"0064682A",
        --14 => X"11A0FFF9",

        ----------------------
        ----- BubbleSort -----
        ----------------------
        --0 => X"34030003",
        --1 => X"AC030000",
        --2 => X"34030004", 
        --3 => X"AC030004",
        --4 => X"34030002",
        --5 => X"AC030008",
        --6 => X"34030001",
        --7 => X"AC03000C",
        --8 => X"34030007",
        --9 => X"AC030010",

        --10 => X"34090014",
        --11 => X"34020000",
        --12 => X"34030000",

        --13 => X"8C440000",
        --14 => X"8C650000",
        --15 => X"0085302A",
        --16 => X"10C00002",
        --17 => X"AC640000",
        --18 => X"AC450000",

        --19 => X"20420004",
        --20 => X"1449FFF8",

        --21 => X"20630004",
        --22 => X"34620000",
        --23 => X"1469FFF5",

        --24 => X"8C070000",
        --25 => X"8C070004",
        --26 => X"8C070008",
        --27 => X"8C07000C",
        --28 => X"8C070010",

        ----------------------
        ----- BinarySort -----
        ----------------------
        --0 => X"34030003",
        --1 => X"AC030000",
        --2 => X"34030004", 
        --3 => X"AC030004",
        --4 => X"34030002",
        --5 => X"AC030008",
        --6 => X"34030001",
        --7 => X"AC03000C",
        --8 => X"34030007",
        --9 => X"AC030010",

        --10 => X"34090014",
        --11 => X"34020000",
        --12 => X"34030000",

        --13 => X"8C440000",
        --14 => X"8C450004",
        --15 => X"0085302A",
        --16 => X"14C00002",
        --17 => X"AC440004",
        --18 => X"AC450000",

        --19 => X"20420004",
        --20 => X"1449FFF8",

        --21 => X"20630004",
        --22 => X"34020000",
        --23 => X"1469FFF5",

        --24 => X"8C070000",
        --25 => X"8C070004",
        --26 => X"8C070008",
        --27 => X"8C07000C",
        --28 => X"8C070010",
        --29 => X"8C070014",


        ----------------------
        -- Bubblesort(mult) --
        ----------------------
        --0 => X"34030003",
        --1 => X"AC030000",
        --2 => X"34030004",
        --3 => X"AC030004",
        --4 => X"34030002",
        --5 => X"AC030008",
        --6 => X"34030001",
        --7 => X"AC03000C",
        --8 => X"34030007",
        --9 => X"AC030010",

        --10 => X"34090005",
        --11 => X"340E0004",
        --12 => X"34020000",
        --13 => X"34030000",

        --14 => X"004E0018",
        --15 => X"00007812",
        --16 => X"8DE40000",
        --17 => X"006E0018",
        --18 => X"00007812",
        --19 => X"8DE50000",
        --20 => X"0085302A",
        --21 => X"10C00006",
        --22 => X"006E0018",
        --23 => X"00007812",
        --24 => X"ADE40000",
        --25 => X"004E0018",
        --26 => X"00007812",
        --27 => X"ADE50000",

        --28 => X"20420001",
        --29 => X"1449FFF0",

        --30 => X"20630001",
        --31 => X"34620000",
        --32 => X"1469FFED",

        --33 => X"8C070000",
        --34 => X"8C070004",
        --35 => X"8C070008",
        --36 => X"8C07000C",
        --37 => X"8C070010",

        ----------------------
        ------ Link Reg ------
        ----------------------
        0 => X"20010001",
        1 => X"20220001",
        2 => X"20430001", 
        3 => X"34050003",

        4 => X"04B10002",
        5 => X"0C000009",
        6 => X"08000004",

        7 => X"00A12822",
        8 => X"03E00008",

        9 => X"03E00008",

        ----------------------
        -------- Misc --------
        ----------------------
        --0 => X"20010005",
        --1 => X"AC010000",
        --2 => X"8C020000", 
        --3 => X"AC020004", 
        --4 => X"8C030000",
        --5 => X"AC620003",
        --6 => X"8C070008",

        --0 => X"20020005",
        --1 => X"2001000A",
        --2 => X"2021FFFF", 
        --3 => X"0421FFFE", 
        --4 => X"20210001",
        --5 => X"0041182A",
        --6 => X"1060FFFD",
        --7 => X"AC230003",

        --0 => X"2001001C",
        --1 => X"2002002F",
        --2 => X"00220018", 
        --3 => X"00001812",
        --4 => X"0020F809",
        --5 => X"00412022",
        --6 => X"000228C0",
        --7 => X"03E00008",
        --0 => X"00231022",
        --1 => X"00456024",
        --2 => X"00c26825",
        --3 => X"00427020",
        --4 => X"ac4f0064",
        --5 => X"00220820",
        --6 => X"00230820",
        --7 => X"00240820",
        --8 => X"8c220014",
        --9 => X"00452024",
        --10 => X"00464025",
        --11 => X"00824820",
        --12 => X"00c7082a",

        others => X"00000000"

    );

begin

    process(CLK)
    begin
        if (RISING_EDGE(CLK)) then
            if (WE = '1') then
                imem(CONV_INTEGER(ADDR)) <= DI;
            end if;
            DO <= imem(CONV_INTEGER(ADDR));
        end if;
    end process;

end IMEM_BR512X32_BEH;

